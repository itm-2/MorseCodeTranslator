module lcd_pos_control (
    input wire clk,           // 50MHz System Clock
    input wire rst_n,         // Active Low Reset
    
    // --- ����� �Է� �������̽� ---
    input wire start_btn,     // 1�� �Ǹ� ���� ���� (��ư ����)
    input wire [3:0] in_col,  // ���� ��ǥ (0 ~ 15) -> ����ġ ����
    input wire [0:0] in_row,  // ���� ��ǥ (0: ����, 1: �Ʒ���) -> ����ġ ����
    
    // --- LCD �ϵ���� �� ---
    output reg lcd_rs,
    output reg lcd_rw,
    output reg lcd_e,
    output reg [7:0] lcd_data
);

    // -------------------------------------------------------------------------
    // �Ķ���� �� ��� ���� (50MHz Ŭ�� ����)
    // -------------------------------------------------------------------------
    parameter CLK_FREQ = 50_000_000;
    
    // Ÿ�̹� ���
    localparam CNT_15MS  = 750_000; 
    localparam CNT_5MS   = 250_000; 
    localparam CNT_100US = 5_000;   
    localparam CNT_CMD   = 2_500;   // 50us (��ɾ� ���� �ð�)
    localparam CNT_CLR   = 100_000; // 2ms (Clear ��ɾ� ���� �ð�)

    // ��ɾ� ����
    localparam CMD_WAKEUP     = 8'h30;
    localparam CMD_FUNC_SET   = 8'h38; // 8-bit, 2-line, 5x8 font
    localparam CMD_DISP_OFF   = 8'h08; 
    localparam CMD_DISP_CLEAR = 8'h01; 
    localparam CMD_ENTRY_MODE = 8'h06; // Auto Increment
    localparam CMD_DISP_ON    = 8'h0C; // Display On, Cursor Off

    // ���� �ӽ� ����
    localparam S_PWR_WAIT   = 0;
    localparam S_INIT_1     = 1;
    localparam S_INIT_2     = 2;
    localparam S_INIT_3     = 3;
    localparam S_FUNC_SET   = 4;
    localparam S_DISP_OFF   = 5;
    localparam S_DISP_CLR   = 6;
    localparam S_ENTRY_MODE = 7;
    localparam S_DISP_ON    = 8;
    localparam S_IDLE       = 9;  // �Է� ��� ����
    localparam S_SET_ADDR   = 10; // ��ǥ ����
    localparam S_WRITE_DATA = 11; // "HELLO WORLD" ���
    localparam S_DONE_WAIT  = 12; // ��ư �� ������ ��� (�ߺ� ����)

    reg [4:0] state;
    reg [31:0] wait_cnt;
    reg [3:0] char_idx; 

    // ����� �޽��� ���� ("HELLO WORLD" - 11����)
    reg [7:0] message [0:10];
    
    // ��ǥ ���� ����
    reg [6:0] target_addr;

    initial begin
        message[0] = "H"; message[1] = "E"; message[2] = "L"; message[3] = "L";
        message[4] = "O"; message[5] = " "; message[6] = "W"; message[7] = "O";
        message[8] = "R"; message[9] = "L"; message[10] = "D";
    end

    // -------------------------------------------------------------------------
    // ���� ����
    // -------------------------------------------------------------------------
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= S_PWR_WAIT;
            wait_cnt <= 0;
            char_idx <= 0;
            lcd_e <= 0; lcd_rs <= 0; lcd_rw <= 0; lcd_data <= 0;
        end else begin
            case (state)
                // ============================================================
                // 1. �ʱ�ȭ ������ (���� ���� �� �ڵ� ����)
                // ============================================================
                S_PWR_WAIT: begin
                    if (wait_cnt >= CNT_15MS) begin wait_cnt <= 0; state <= S_INIT_1; end
                    else wait_cnt <= wait_cnt + 1;
                end

                S_INIT_1: begin // 0x30
                    lcd_rs <= 0; lcd_rw <= 0; lcd_data <= CMD_WAKEUP;
                    if (wait_cnt == 2) lcd_e <= 1; else if (wait_cnt == 22) lcd_e <= 0; // Timing Fix
                    if (wait_cnt >= (CNT_5MS + 22)) begin wait_cnt <= 0; state <= S_INIT_2; end
                    else wait_cnt <= wait_cnt + 1;
                end

                S_INIT_2: begin // 0x30
                    lcd_rs <= 0; lcd_rw <= 0; lcd_data <= CMD_WAKEUP;
                    if (wait_cnt == 2) lcd_e <= 1; else if (wait_cnt == 22) lcd_e <= 0;
                    if (wait_cnt >= (CNT_100US + 22)) begin wait_cnt <= 0; state <= S_INIT_3; end
                    else wait_cnt <= wait_cnt + 1;
                end

                S_INIT_3: begin // 0x30
                    lcd_rs <= 0; lcd_rw <= 0; lcd_data <= CMD_WAKEUP;
                    if (wait_cnt == 2) lcd_e <= 1; else if (wait_cnt == 22) lcd_e <= 0;
                    if (wait_cnt >= (CNT_CMD + 22)) begin wait_cnt <= 0; state <= S_FUNC_SET; end
                    else wait_cnt <= wait_cnt + 1;
                end

                S_FUNC_SET: begin // 0x38
                    lcd_rs <= 0; lcd_rw <= 0; lcd_data <= CMD_FUNC_SET;
                    if (wait_cnt == 2) lcd_e <= 1; else if (wait_cnt == 22) lcd_e <= 0;
                    if (wait_cnt >= (CNT_CMD + 22)) begin wait_cnt <= 0; state <= S_DISP_OFF; end
                    else wait_cnt <= wait_cnt + 1;
                end

                S_DISP_OFF: begin // 0x08
                    lcd_rs <= 0; lcd_rw <= 0; lcd_data <= CMD_DISP_OFF;
                    if (wait_cnt == 2) lcd_e <= 1; else if (wait_cnt == 22) lcd_e <= 0;
                    if (wait_cnt >= (CNT_CMD + 22)) begin wait_cnt <= 0; state <= S_DISP_CLR; end
                    else wait_cnt <= wait_cnt + 1;
                end

                S_DISP_CLR: begin // 0x01
                    lcd_rs <= 0; lcd_rw <= 0; lcd_data <= CMD_DISP_CLEAR;
                    if (wait_cnt == 2) lcd_e <= 1; else if (wait_cnt == 22) lcd_e <= 0;
                    if (wait_cnt >= (CNT_CLR + 22)) begin wait_cnt <= 0; state <= S_ENTRY_MODE; end
                    else wait_cnt <= wait_cnt + 1;
                end

                S_ENTRY_MODE: begin // 0x06
                    lcd_rs <= 0; lcd_rw <= 0; lcd_data <= CMD_ENTRY_MODE;
                    if (wait_cnt == 2) lcd_e <= 1; else if (wait_cnt == 22) lcd_e <= 0;
                    if (wait_cnt >= (CNT_CMD + 22)) begin wait_cnt <= 0; state <= S_DISP_ON; end
                    else wait_cnt <= wait_cnt + 1;
                end

                S_DISP_ON: begin // 0x0C
                    lcd_rs <= 0; lcd_rw <= 0; lcd_data <= CMD_DISP_ON;
                    if (wait_cnt == 2) lcd_e <= 1; else if (wait_cnt == 22) lcd_e <= 0;
                    if (wait_cnt >= (CNT_CMD + 22)) begin wait_cnt <= 0; state <= S_IDLE; end
                    else wait_cnt <= wait_cnt + 1;
                end

                // ============================================================
                // 2. ��� �� ����� �Է� ó��
                // ============================================================
                S_IDLE: begin
                    lcd_e <= 0;
                    wait_cnt <= 0;
                    
                    // ��ư�� ������ ��ǥ ��� �� �̵� ����
                    if (start_btn == 1'b1) begin
                        // [��ǥ ��� ����]
                        // Row 0: 0x00 ~ 0x0F
                        // Row 1: 0x40 ~ 0x4F
                        if (in_row == 1'b0) target_addr <= {3'b000, in_col}; // 0x00 + col
                        else                target_addr <= {3'b100, in_col}; // 0x40 + col
                        
                        state <= S_SET_ADDR;
                    end
                end

                // 3. Ŀ�� ��ġ ���� (Set DDRAM Address)
                S_SET_ADDR: begin
                    lcd_rs <= 0; lcd_rw <= 0;
                    lcd_data <= {1'b1, target_addr}; // Command: 0x80 | Address

                    if (wait_cnt == 2) lcd_e <= 1; else if (wait_cnt == 22) lcd_e <= 0;

                    if (wait_cnt >= (CNT_CMD + 22)) begin
                        wait_cnt <= 0;
                        char_idx <= 0;
                        state <= S_WRITE_DATA;
                    end else wait_cnt <= wait_cnt + 1;
                end

                // 4. "HELLO WORLD" ��� ����
                S_WRITE_DATA: begin
                    lcd_rs <= 1; // Data ���
                    lcd_rw <= 0;
                    lcd_data <= message[char_idx];

                    if (wait_cnt == 2) lcd_e <= 1; else if (wait_cnt == 22) lcd_e <= 0;

                    if (wait_cnt >= (CNT_CMD + 22)) begin
                        wait_cnt <= 0;
                        // 11���� (0~10) �� ������ ����
                        if (char_idx == 10) state <= S_DONE_WAIT;
                        else char_idx <= char_idx + 1;
                    end else wait_cnt <= wait_cnt + 1;
                end

                // 5. ��ư �� ������ ��� (�ߺ� ���� ����)
                S_DONE_WAIT: begin
                    lcd_e <= 0;
                    if (start_btn == 1'b0) begin
                        state <= S_IDLE; // ��ư�� ���� �ٽ� �Է� ��� ���·�
                    end
                end

                default: state <= S_PWR_WAIT;
            endcase
        end
    end

endmodule