`timescale 1ns / 1ps

module tb_MorseSystem_Fast;

    // Ŭ�� & ����
    reg clk;
    reg rst_n;
    
    // �Է� ��ȣ�� - �ʱⰪ ���!
    reg [4:0] btn = 5'b00000;           // �� �ʱⰪ �߰�
    reg [2:0] speed_sel = 3'b000;       // �� �ʱⰪ �߰�
    reg is_active = 1'b0;               // �� �ʱⰪ �߰�
    
    // ��� ��ȣ��
    wire [9:0] led;
    wire [2:0] rgb_r, rgb_g, rgb_b;
    wire piezo;
    wire servo;
    wire lcd_e, lcd_rs, lcd_rw;
    wire [7:0] lcd_data;

    // DUT �ν��Ͻ�
    MorseSystemTop #(
        .CLK_HZ(100_000_000)
    ) dut (
        .clk(clk),
        .rst_n(rst_n),
        .btn(btn),
        .speed_sel(speed_sel),
        .is_active(is_active),
        .led(led),
        .rgb_r(rgb_r),
        .rgb_g(rgb_g),
        .rgb_b(rgb_b),
        .piezo(piezo),
        .servo(servo),
        .lcd_e(lcd_e),
        .lcd_rs(lcd_rs),
        .lcd_rw(lcd_rw),
        .lcd_data(lcd_data)
    );

    // Ŭ�� ���� (100MHz = 10ns)
    initial begin
        clk = 0;  // �� ����� �ʱ�ȭ
        forever #5 clk = ~clk;
    end

    // ���� ������ ��ȭ
    initial begin
        // �ʱ� ����
        rst_n = 0;
        btn = 5'b00000;
        speed_sel = 3'b000;
        is_active = 0;
        
        // ����� ���� �ð�
        #200;
        
        // ���� ����
        rst_n = 1;
        #100;
        
        // �ý��� Ȱ��ȭ
        is_active = 1;
        #100;
        
        $display("=== Initialization Complete ===");
        $display("Time: %0t", $time);
        $display("rst_n: %b", rst_n);
        $display("is_active: %b", is_active);
        $display("LED: %b", led);
        
        // ������ �׽�Ʈ
        $display("\n=== Button Test ===");
        btn = 5'b00001;
        #100;
        btn = 5'b00000;
        #100;
        
        $display("Test complete!");
        $finish;
    end

    // Ÿ�Ӿƿ�
    initial begin
        #10000;
        $display("Timeout!");
        $finish;
    end

    // ��ȣ ����͸�
    initial begin
        $monitor("Time=%0t rst_n=%b btn=%b led=%b", 
                 $time, rst_n, btn, led);
    end

endmodule