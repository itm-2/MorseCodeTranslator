module morse_decoder_final (
    input wire clk,           // 50MHz System Clock
    input wire rst_n,         // Active Low Reset
    
    // --- Input Keys ---
    input wire btn_key,       // �� ��ȣ �Է� Ű (Morse Input)
    input wire btn_enter,     // ��� Ȯ�� / ��� ��ȯ
    input wire btn_back,      // �ڷ� ����
    input wire btn_up,        // ������ �� (Result ȭ���)
    input wire btn_down,      // ������ �ٿ� (Result ȭ���)

    // --- Output ---
    output reg [3:0] led,     // LED ��� (WarnInvalid, KeyFeedback)
    
    // --- LCD Interface ---
    output wire lcd_rs,
    output wire lcd_rw,
    output wire lcd_e,
    output wire [7:0] lcd_data
);

    // =========================================================================
    // 1. �Ķ���� �� ��� ���� (UserSetting �ݿ�)
    // =========================================================================
    parameter CLK_FREQ = 50_000_000;
    
    // KeyMapping & Action Settings
    // 1ms = 50,000 clk
    localparam THRESHOLD_DIT_DAH = 10_000_000; // 200ms (����: Dit, �ʰ�: Dah)
    localparam THRESHOLD_GAP     = 25_000_000; // 500ms (���� ���� Space ����)
    
    // UI ���� ���� (UUID ���� ��ü)
    localparam S_INTRO      = 0; // "ENTER THE CODE..."
    localparam S_DECODE     = 1; // �ǽð� �Է� �� �ص�
    localparam S_RESULT     = 2; // ��ü ��� ��ȸ (Paging)
    
    // =========================================================================
    // 2. ���� ���� �� ��������
    // =========================================================================
    reg [2:0]  ui_state;      // ���� UI ����
    
    // Ÿ�̸� �� Ű ó��
    reg [31:0] timer_press;   // KeyAction: ���� �ð�
    reg [31:0] timer_gap;     // KeyAction: �� �ð� (AutoDitGap)
    reg key_prev;             // Edge Detection��
    
    // �� ��ȣ ���� ���� (IBuffer ����)
    // �ִ� 6���� ��ȣ (����/Ư������ ����) ����. 0:Dit, 1:Dah
    reg [5:0] pattern_reg;    
    reg [2:0] pattern_len;    
    
    // �ؽ�Ʈ ���� (Buffer ����) - �ִ� 128���� ����
    reg [7:0] text_buffer [0:127]; 
    reg [6:0] buf_head;       // ���� ���� ��ġ
    reg [6:0] page_idx;       // ��� ȭ�� ����¡ �ε���

    // LCD ǥ�ÿ� ���� ����
    reg [127:0] lcd_line1;
    reg [127:0] lcd_line2;

    // WarnInvalid (LED ����)
    reg [31:0] warn_timer;
    reg is_warning;

    // ��ư Debounce �� One-shot ó���� ���� ��������
    reg btn_enter_prev, btn_back_prev, btn_up_prev, btn_down_prev;
    
    // =========================================================================
    // 3. ���� ���� (Always Block)
    // =========================================================================
    
    // Translator Function (���� ��)
    function [7:0] translate_morse;
        input [2:0] len;
        input [5:0] pat; // LSB�� ù �Է� (Shift��)
        begin
            case ({len, pat})
                // Length 1
                {3'd1, 6'b00000_0}: translate_morse = "E"; // .
                {3'd1, 6'b00000_1}: translate_morse = "T"; // -
                // Length 2
                {3'd2, 6'b0000_01}: translate_morse = "A"; // .-
                {3'd2, 6'b0000_10}: translate_morse = "N"; // -.
                {3'd2, 6'b0000_00}: translate_morse = "I"; // ..
                {3'd2, 6'b0000_11}: translate_morse = "M"; // --
                // Length 3
                {3'd3, 6'b000_000}: translate_morse = "S"; // ...
                {3'd3, 6'b000_111}: translate_morse = "O"; // ---
                {3'd3, 6'b000_010}: translate_morse = "R"; // .-.
                {3'd3, 6'b000_100}: translate_morse = "D"; // -..
                {3'd3, 6'b000_101}: translate_morse = "K"; // -.-
                {3'd3, 6'b000_110}: translate_morse = "G"; // --.
                {3'd3, 6'b000_001}: translate_morse = "U"; // ..-
                {3'd3, 6'b000_011}: translate_morse = "W"; // .--
                // Length 4 (���� �Ϻ�)
                {3'd4, 6'b00_0000}: translate_morse = "H"; // ....
                {3'd4, 6'b00_1010}: translate_morse = "C"; // -.-.
                {3'd4, 6'b00_0111}: translate_morse = "J"; // .---
                {3'd4, 6'b00_1101}: translate_morse = "Q"; // --.-
                {3'd4, 6'b00_1011}: translate_morse = "Y"; // -.--
                {3'd4, 6'b00_0001}: translate_morse = "V"; // ...-
                {3'd4, 6'b00_1000}: translate_morse = "B"; // -...
                {3'd4, 6'b00_0100}: translate_morse = "L"; // .-..
                {3'd4, 6'b00_0010}: translate_morse = "F"; // ..-.
                {3'd4, 6'b00_0101}: translate_morse = "+"; // .-.- (AR)
                default: translate_morse = 0; // Invalid
            endcase
        end
    endfunction

    reg [7:0] decoded_char; // ���� ��� �ӽ� ����

    integer i;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            ui_state <= S_INTRO;
            timer_press <= 0; timer_gap <= 0;
            key_prev <= 0;
            pattern_reg <= 0; pattern_len <= 0;
            buf_head <= 0; page_idx <= 0;
            is_warning <= 0; warn_timer <= 0;
            // ���� �ʱ�ȭ (�ռ� �ÿ� ���õ� �� ����, ���ۻ� ����� �ϹǷ� ����)
            for(i=0; i<128; i=i+1) text_buffer[i] <= " "; 
        end else begin
            // Edge Detection
            btn_enter_prev <= btn_enter;
            btn_back_prev <= btn_back;
            btn_up_prev <= btn_up;
            btn_down_prev <= btn_down;
            key_prev <= btn_key;

            // --- WarnInvalid Timer ---
            if (is_warning) begin
                if (warn_timer > 0) warn_timer <= warn_timer - 1;
                else is_warning <= 0;
            end

            // --- UI State Machine ---
            case (ui_state)
                // ------------------------------------------------------------
                // [ȭ�� 0] �ʱ� ȭ��: "ENTER THE CODE..."
                // ------------------------------------------------------------
                S_INTRO: begin
                    if (btn_key || (btn_enter && !btn_enter_prev)) begin
                        // �ƹ� Ű�� ������ ���ڵ� ȭ������ ��ȯ
                        ui_state <= S_DECODE;
                        buf_head <= 0;
                        pattern_len <= 0;
                        pattern_reg <= 0;
                        // ���� Clear
                        for(i=0; i<128; i=i+1) text_buffer[i] <= " ";
                    end
                end

                // ------------------------------------------------------------
                // [ȭ�� 1] Decoding: �ǽð� �Է� �� �ص�
                // ------------------------------------------------------------
                S_DECODE: begin
                    // 1. KeyAction Logic (Dit/Dah Detection)
                    if (btn_key) begin // ������ ���� ��
                        timer_press <= timer_press + 1;
                        timer_gap <= 0; // �� Ÿ�̸� ����
                    end else begin // ���� ���� ��
                        // Falling Edge ���� (��ư �� ����)
                        if (key_prev == 1'b1) begin
                            if (timer_press > THRESHOLD_DIT_DAH) begin
                                // Dah (10 -> 1�� ����)
                                pattern_reg <= {pattern_reg[4:0], 1'b1}; 
                            end else begin
                                // Dit (01 -> 0���� ����)
                                pattern_reg <= {pattern_reg[4:0], 1'b0};
                            end
                            pattern_len <= pattern_len + 1;
                            timer_press <= 0;
                        end

                        // Gap Detection (Space ����)
                        if (pattern_len > 0) begin
                            timer_gap <= timer_gap + 1;
                            
                            // UserSetting�� DitGap��ŭ ��� �� ����
                            if (timer_gap > THRESHOLD_GAP) begin
                                // Translator ȣ��
                                decoded_char = translate_morse(pattern_len, pattern_reg);
                                
                                if (decoded_char != 0) begin
                                    // ��ȿ�� ���� -> Buffer Push
                                    text_buffer[buf_head] <= decoded_char;
                                    buf_head <= buf_head + 1;
                                end else begin
                                    // Invalid (0 ��ȯ��) -> warnInvalid
                                    is_warning <= 1;
                                    warn_timer <= CLK_FREQ / 2; // 0.5��
                                end
                                
                                // �� ���� �ʱ�ȭ
                                pattern_reg <= 0;
                                pattern_len <= 0;
                                timer_gap <= 0;
                            end
                        end
                    end

                    // 2. Navigation
                    if (btn_enter && !btn_enter_prev) begin
                        ui_state <= S_RESULT;
                        page_idx <= 0; // ù ����������
                    end
                    if (btn_back && !btn_back_prev) begin
                        ui_state <= S_INTRO;
                    end
                end

                // ------------------------------------------------------------
                // [ȭ�� 2] Result: ��ü ��� Ȯ�� (Paging)
                // ------------------------------------------------------------
                S_RESULT: begin
                    // Navigation
                    if (btn_enter && !btn_enter_prev) begin
                        ui_state <= S_DECODE; // �ٽ� ���ڵ� ȭ������
                    end
                    if (btn_back && !btn_back_prev) begin
                        ui_state <= S_DECODE; // ���� ȭ������
                    end

                    // Paging (UP/DOWN) - 15���� ����
                    if (btn_down && !btn_down_prev) begin
                        if (page_idx + 15 < buf_head) 
                            page_idx <= page_idx + 15;
                    end
                    if (btn_up && !btn_up_prev) begin
                        if (page_idx >= 15)
                            page_idx <= page_idx - 15;
                        else
                            page_idx <= 0;
                    end
                end
            endcase
        end
    end

    // =========================================================================
    // 4. Output Logic (LED & LCD)
    // =========================================================================

    // LED: printLED (KeyMap) + warnInvalid
    always @(*) begin
        if (is_warning) begin
            led = 4'b1111; // ��� �� ��ü ����
        end else begin
            // printLED: ��� ������ ��ư ��Ī
            // ��: Intro���� Enter��, Decode���� Key/Enter/Back ��
            case (ui_state)
                S_INTRO:  led = {btn_key, 3'b000}; 
                S_DECODE: led = {btn_key, 1'b0, 1'b0, 1'b0}; // �Է� �� ����
                S_RESULT: led = 4'b0000; // ��� ȭ�鿡�� �ҵ�
                default:  led = 4'b0000;
            endcase
        end
    end

    // LCD Buffer Mapping (showUI)
    always @(*) begin
        // �⺻�� ���� ä��
        lcd_line1 = {16{8'h20}};
        lcd_line2 = {16{8'h20}};

        case (ui_state)
            S_INTRO: begin
                lcd_line1 = "ENTER THE CODE.."; // �߾� ���� ����
                lcd_line2 = "PRESS ANY KEY   ";
            end

            S_DECODE: begin
                // Row 1: ������� �Էµ� �ؽ�Ʈ�� ���κ� (�ֱ� 16��)
                // 15���� ������ �� 0����, �Ѿ�� ��ũ��
                for (i=0; i<16; i=i+1) begin
                    if (buf_head < 16) begin
                        if (i < buf_head) lcd_line1[127 - i*8 -: 8] = text_buffer[i];
                    end else begin
                        // ������ 16���� �����ֱ�
                        lcd_line1[127 - i*8 -: 8] = text_buffer[buf_head - 16 + i];
                    end
                end

                // Row 2: ���� �Է� ���� �� ��ȣ ���� (.-...)
                for (i=0; i<6; i=i+1) begin
                    if (i < pattern_len) begin
                        // LSB���� �ԷµǾ����Ƿ� ���� ���� (���⼱ ���ǻ� 0���� ���)
                        if (pattern_reg[pattern_len - 1 - i] == 1) 
                             lcd_line2[127 - i*8 -: 8] = "-"; // Dah
                        else lcd_line2[127 - i*8 -: 8] = "."; // Dit
                    end
                end
            end

            S_RESULT: begin
                // Row 1: page_idx ���� 15����
                // Row 2: page_idx+15 ���� 15���� (prompt: "Buffer�� page ����(15����)")
                for (i=0; i<16; i=i+1) begin
                    // Line 1
                    if (page_idx + i < 128)
                        lcd_line1[127 - i*8 -: 8] = text_buffer[page_idx + i];
                    
                    // Line 2 (���� ������ �̸����� ���� Ȥ�� ���� ���)
                    if (page_idx + 15 + i < 128)
                        lcd_line2[127 - i*8 -: 8] = text_buffer[page_idx + 15 + i];
                end
            end
        endcase
    end

    // LCD Driver �ν��Ͻ�
    lcd_driver_ctrl u_lcd (
        .clk(clk),
        .rst_n(rst_n),
        .line1(lcd_line1),
        .line2(lcd_line2),
        .lcd_rs(lcd_rs),
        .lcd_rw(lcd_rw),
        .lcd_e(lcd_e),
        .lcd_data(lcd_data)
    );

endmodule


// =============================================================================
// LCD Driver Module (������Ʈ�� ������ ���� ���)
// =============================================================================
module lcd_driver_ctrl (
    input wire clk,
    input wire rst_n,
    input wire [127:0] line1,
    input wire [127:0] line2,
    output reg lcd_rs,
    output reg lcd_rw,
    output reg lcd_e,
    output reg [7:0] lcd_data
);
    // Ÿ�̹� �Ķ���� (50MHz)
    localparam CNT_CMD = 2_500;   
    localparam CNT_INIT_WAIT = 2_000_000; // 40ms

    reg [3:0] state;
    reg [31:0] cnt;
    reg [3:0] char_idx; 
    reg line_sel;       

    localparam S_INIT_PWR  = 0;
    localparam S_FUNC_SET  = 1;
    localparam S_DISP_ON   = 2;
    localparam S_CLR       = 3;
    localparam S_MODE      = 4;
    localparam S_ADDR      = 5;
    localparam S_WRITE     = 6;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= S_INIT_PWR;
            cnt <= 0; char_idx <= 0; line_sel <= 0;
            lcd_e <= 0; lcd_rs <= 0; lcd_rw <= 0;
        end else begin
            case (state)
                S_INIT_PWR: begin // Power Wait
                    if (cnt > CNT_INIT_WAIT) begin cnt <= 0; state <= S_FUNC_SET; end
                    else cnt <= cnt + 1;
                end
                S_FUNC_SET: begin // 0x38
                    lcd_rs <= 0; lcd_rw <= 0; lcd_data <= 8'h38;
                    if (cnt == 2) lcd_e <= 1; else if (cnt == 22) lcd_e <= 0;
                    if (cnt > CNT_CMD + 22) begin cnt <= 0; state <= S_DISP_ON; end
                    else cnt <= cnt + 1;
                end
                S_DISP_ON: begin // 0x0C
                    lcd_rs <= 0; lcd_rw <= 0; lcd_data <= 8'h0C;
                    if (cnt == 2) lcd_e <= 1; else if (cnt == 22) lcd_e <= 0;
                    if (cnt > CNT_CMD + 22) begin cnt <= 0; state <= S_CLR; end
                    else cnt <= cnt + 1;
                end
                S_CLR: begin // 0x01
                    lcd_rs <= 0; lcd_rw <= 0; lcd_data <= 8'h01;
                    if (cnt == 2) lcd_e <= 1; else if (cnt == 22) lcd_e <= 0;
                    if (cnt > 100_000 + 22) begin cnt <= 0; state <= S_MODE; end // Clear is slow
                    else cnt <= cnt + 1;
                end
                S_MODE: begin // 0x06
                    lcd_rs <= 0; lcd_rw <= 0; lcd_data <= 8'h06;
                    if (cnt == 2) lcd_e <= 1; else if (cnt == 22) lcd_e <= 0;
                    if (cnt > CNT_CMD + 22) begin cnt <= 0; state <= S_ADDR; end
                    else cnt <= cnt + 1;
                end

                // --- Refresh Loop ---
                S_ADDR: begin
                    lcd_rs <= 0; lcd_rw <= 0;
                    if (line_sel == 0) lcd_data <= 8'h80 + char_idx; // Line 1
                    else               lcd_data <= 8'hC0 + char_idx; // Line 2

                    if (cnt == 2) lcd_e <= 1; else if (cnt == 22) lcd_e <= 0;
                    if (cnt > CNT_CMD + 22) begin cnt <= 0; state <= S_WRITE; end
                    else cnt <= cnt + 1;
                end
                S_WRITE: begin
                    lcd_rs <= 1; lcd_rw <= 0;
                    if (line_sel == 0) lcd_data <= line1[127 - char_idx*8 -: 8];
                    else               lcd_data <= line2[127 - char_idx*8 -: 8];

                    if (cnt == 2) lcd_e <= 1; else if (cnt == 22) lcd_e <= 0;
                    if (cnt > CNT_CMD + 22) begin 
                        cnt <= 0;
                        if (char_idx == 15) begin
                            char_idx <= 0;
                            line_sel <= ~line_sel; // �� �ٲ�
                        end else begin
                            char_idx <= char_idx + 1;
                        end
                        state <= S_ADDR;
                    end else cnt <= cnt + 1;
                end
            endcase
        end
    end
endmodule